`timescale 1ns / 1ps

module alpha(
    input [31:0] alpha_in,
    output [31:0] alpha_out
    );
    wire [31:0] lut_out;
    wire [31:0] shift_out;
    
    reg [8:0] t0=8'd0;
    reg [8:0] t1=8'd0;
    reg [8:0] t2=8'd0;
    reg [8:0] t3=8'd0;
  
    function [7 : 0] al(input [7 : 0] z);
    begin
      case (z)
        8'h00: al = 8'h63;
        8'h01: al = 8'h7c;
        8'h02: al = 8'h77;
        8'h03: al = 8'h7b;
        8'h04: al = 8'hf2;
        8'h05: al = 8'h6b;
        8'h06: al = 8'h6f;
        8'h07: al = 8'hc5;
        8'h08: al = 8'h30;
        8'h09: al = 8'h01;
        8'h0a: al = 8'h67;
        8'h0b: al = 8'h2b;
        8'h0c: al = 8'hfe;
        8'h0d: al = 8'hd7;
        8'h0e: al = 8'hab;
        8'h0f: al = 8'h76;
        8'h10: al = 8'hca;
        8'h11: al = 8'h82;
        8'h12: al = 8'hc9;
        8'h13: al = 8'h7d;
        8'h14: al = 8'hfa;
        8'h15: al = 8'h59;
        8'h16: al = 8'h47;
        8'h17: al = 8'hf0;
        8'h18: al = 8'had;
        8'h19: al = 8'hd4;
        8'h1a: al = 8'ha2;
        8'h1b: al = 8'haf;
        8'h1c: al = 8'h9c;
        8'h1d: al = 8'ha4;
        8'h1e: al = 8'h72;
        8'h1f: al = 8'hc0;
        8'h20: al = 8'hb7;
        8'h21: al = 8'hfd;
        8'h22: al = 8'h93;
        8'h23: al = 8'h26;
        8'h24: al = 8'h36;
        8'h25: al = 8'h3f;
        8'h26: al = 8'hf7;
        8'h27: al = 8'hcc;
        8'h28: al = 8'h34;
        8'h29: al = 8'ha5;
        8'h2a: al = 8'he5;
        8'h2b: al = 8'hf1;
        8'h2c: al = 8'h71;
        8'h2d: al = 8'hd8;
        8'h2e: al = 8'h31;
        8'h2f: al = 8'h15;
        8'h30: al = 8'h04;
        8'h31: al = 8'hc7;
        8'h32: al = 8'h23;
        8'h33: al = 8'hc3;
        8'h34: al = 8'h18;
        8'h35: al = 8'h96;
        8'h36: al = 8'h05;
        8'h37: al = 8'h9a;
        8'h38: al = 8'h07;
        8'h39: al = 8'h12;
        8'h3a: al = 8'h80;
        8'h3b: al = 8'he2;
        8'h3c: al = 8'heb;
        8'h3d: al = 8'h27;
        8'h3e: al = 8'hb2;
        8'h3f: al = 8'h75;
        8'h40: al = 8'h09;
        8'h41: al = 8'h83;
        8'h42: al = 8'h2c;
        8'h43: al = 8'h1a;
        8'h44: al = 8'h1b;
        8'h45: al = 8'h6e;
        8'h46: al = 8'h5a;
        8'h47: al = 8'ha0;
        8'h48: al = 8'h52;
        8'h49: al = 8'h3b;
        8'h4a: al = 8'hd6;
        8'h4b: al = 8'hb3;
        8'h4c: al = 8'h29;
        8'h4d: al = 8'he3;
        8'h4e: al = 8'h2f;
        8'h4f: al = 8'h84;
        8'h50: al = 8'h53;
        8'h51: al = 8'hd1;
        8'h52: al = 8'h00;
        8'h53: al = 8'hed;
        8'h54: al = 8'h20;
        8'h55: al = 8'hfc;
        8'h56: al = 8'hb1;
        8'h57: al = 8'h5b;
        8'h58: al = 8'h6a;
        8'h59: al = 8'hcb;
        8'h5a: al = 8'hbe;
        8'h5b: al = 8'h39;
        8'h5c: al = 8'h4a;
        8'h5d: al = 8'h4c;
        8'h5e: al = 8'h58;
        8'h5f: al = 8'hcf;
        8'h60: al = 8'hd0;
        8'h61: al = 8'hef;
        8'h62: al = 8'haa;
        8'h63: al = 8'hfb;
        8'h64: al = 8'h43;
        8'h65: al = 8'h4d;
        8'h66: al = 8'h33;
        8'h67: al = 8'h85;
        8'h68: al = 8'h45;
        8'h69: al = 8'hf9;
        8'h6a: al = 8'h02;
        8'h6b: al = 8'h7f;
        8'h6c: al = 8'h50;
        8'h6d: al = 8'h3c;
        8'h6e: al = 8'h9f;
        8'h6f: al = 8'ha8;
        8'h70: al = 8'h51;
        8'h71: al = 8'ha3;
        8'h72: al = 8'h40;
        8'h73: al = 8'h8f;
        8'h74: al = 8'h92;
        8'h75: al = 8'h9d;
        8'h76: al = 8'h38;
        8'h77: al = 8'hf5;
        8'h78: al = 8'hbc;
        8'h79: al = 8'hb6;
        8'h7a: al = 8'hda;
        8'h7b: al = 8'h21;
        8'h7c: al = 8'h10;
        8'h7d: al = 8'hff;
        8'h7e: al = 8'hf3;
        8'h7f: al = 8'hd2;
        8'h80: al = 8'hcd;
        8'h81: al = 8'h0c;
        8'h82: al = 8'h13;
        8'h83: al = 8'hec;
        8'h84: al = 8'h5f;
        8'h85: al = 8'h97;
        8'h86: al = 8'h44;
        8'h87: al = 8'h17;
        8'h88: al = 8'hc4;
        8'h89: al = 8'ha7;
        8'h8a: al = 8'h7e;
        8'h8b: al = 8'h3d;
        8'h8c: al = 8'h64;
        8'h8d: al = 8'h5d;
        8'h8e: al = 8'h19;
        8'h8f: al = 8'h73;
        8'h90: al = 8'h60;
        8'h91: al = 8'h81;
        8'h92: al = 8'h4f;
        8'h93: al = 8'hdc;
        8'h94: al = 8'h22;
        8'h95: al = 8'h2a;
        8'h96: al = 8'h90;
        8'h97: al = 8'h88;
        8'h98: al = 8'h46;
        8'h99: al = 8'hee;
        8'h9a: al = 8'hb8;
        8'h9b: al = 8'h14;
        8'h9c: al = 8'hde;
        8'h9d: al = 8'h5e;
        8'h9e: al = 8'h0b;
        8'h9f: al = 8'hdb;
        8'ha0: al = 8'he0;
        8'ha1: al = 8'h32;
        8'ha2: al = 8'h3a;
        8'ha3: al = 8'h0a;
        8'ha4: al = 8'h49;
        8'ha5: al = 8'h06;
        8'ha6: al = 8'h24;
        8'ha7: al = 8'h5c;
        8'ha8: al = 8'hc2;
        8'ha9: al = 8'hd3;
        8'haa: al = 8'hac;
        8'hab: al = 8'h62;
        8'hac: al = 8'h91;
        8'had: al = 8'h95;
        8'hae: al = 8'he4;
        8'haf: al = 8'h79;
        8'hb0: al = 8'he7;
        8'hb1: al = 8'hc8;
        8'hb2: al = 8'h37;
        8'hb3: al = 8'h6d;
        8'hb4: al = 8'h8d;
        8'hb5: al = 8'hd5;
        8'hb6: al = 8'h4e;
        8'hb7: al = 8'ha9;
        8'hb8: al = 8'h6c;
        8'hb9: al = 8'h56;
        8'hba: al = 8'hf4;
        8'hbb: al = 8'hea;
        8'hbc: al = 8'h65;
        8'hbd: al = 8'h7a;
        8'hbe: al = 8'hae;
        8'hbf: al = 8'h08;
        8'hc0: al = 8'hba;
        8'hc1: al = 8'h78;
        8'hc2: al = 8'h25;
        8'hc3: al = 8'h2e;
        8'hc4: al = 8'h1c;
        8'hc5: al = 8'ha6;
        8'hc6: al = 8'hb4;
        8'hc7: al = 8'hc6;
        8'hc8: al = 8'he8;
        8'hc9: al = 8'hdd;
        8'hca: al = 8'h74;
        8'hcb: al = 8'h1f;
        8'hcc: al = 8'h4b;
        8'hcd: al = 8'hbd;
        8'hce: al = 8'h8b;
        8'hcf: al = 8'h8a;
        8'hd0: al = 8'h70;
        8'hd1: al = 8'h3e;
        8'hd2: al = 8'hb5;
        8'hd3: al = 8'h66;
        8'hd4: al = 8'h48;
        8'hd5: al = 8'h03;
        8'hd6: al = 8'hf6;
        8'hd7: al = 8'h0e;
        8'hd8: al = 8'h61;
        8'hd9: al = 8'h35;
        8'hda: al = 8'h57;
        8'hdb: al = 8'hb9;
        8'hdc: al = 8'h86;
        8'hdd: al = 8'hc1;
        8'hde: al = 8'h1d;
        8'hdf: al = 8'h9e;
        8'he0: al = 8'he1;
        8'he1: al = 8'hf8;
        8'he2: al = 8'h98;
        8'he3: al = 8'h11;
        8'he4: al = 8'h69;
        8'he5: al = 8'hd9;
        8'he6: al = 8'h8e;
        8'he7: al = 8'h94;
        8'he8: al = 8'h9b;
        8'he9: al = 8'h1e;
        8'hea: al = 8'h87;
        8'heb: al = 8'he9;
        8'hec: al = 8'hce;
        8'hed: al = 8'h55;
        8'hee: al = 8'h28;
        8'hef: al = 8'hdf;
        8'hf0: al = 8'h8c;
        8'hf1: al = 8'ha1;
        8'hf2: al = 8'h89;
        8'hf3: al = 8'h0d;
        8'hf4: al = 8'hbf;
        8'hf5: al = 8'he6;
        8'hf6: al = 8'h42;
        8'hf7: al = 8'h68;
        8'hf8: al = 8'h41;
        8'hf9: al = 8'h99;
        8'hfa: al = 8'h2d;
        8'hfb: al = 8'h0f;
        8'hfc: al = 8'hb0;
        8'hfd: al = 8'h54;
        8'hfe: al = 8'hbb;
        8'hff: al = 8'h16;
      endcase
    end
    endfunction    
    
    always@(*)
    begin
        t0 <= alpha_in[7:0];
        t1 <= alpha_in[15:8];
        t2 <= alpha_in[23:16];
        t3 <= alpha_in[31:24];
    end
    
    assign shift_out = alpha_in >> 8;
    assign lut_out[7:0] = al(t0);
    assign lut_out[15:8] = al(t1);
    assign lut_out[23:16] = al(t2);
    assign lut_out[31:24] = al(t3);
    assign alpha_out = (lut_out ^ shift_out);
    
endmodule